module main
import hello

fn main() {
    println(hello.hello())
}
