module hello

pub fn hello() string {
    return 'Hello world !'
}

/*
fn main() {
    println(hello())
}
*/
